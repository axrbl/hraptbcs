interface module_common (
    input wire clk,
    input wire rst ;
    ;
    in
    
endinterface //mod